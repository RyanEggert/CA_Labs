// fsm.t.v

module testFSM();
	
endmodule
